
// control unit test bench

module register_module (save,reset,alu_out,data_out);
  reg save;
  reg reset;
  reg [7:0] alu_out;
  wire  [7:0] data_out;
  wire  [7:0] data_out;

  register_module  uut(save,reset,alu_out,data_out);
      initial
           begin
            
           end
endmodule





